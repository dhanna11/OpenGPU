-- OpenGPU Testbench --

entity ogpu_testbench is
end ogpu_testbench;

architecture ogpu_raster_unit_tb1 of ogpu_testbench is
begin
end ogpu_raster_unit_tb1;